library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 
package instructions_core_3 is 
 constant LDA_IMM : std_logic_vector (7 downto 0) :=x"2f"; 
 constant LDB_IMM : std_logic_vector (7 downto 0) :=x"41"; 
 constant LDA_DIR : std_logic_vector (7 downto 0) :=x"a7"; 
 constant LDB_DIR : std_logic_vector (7 downto 0) :=x"12"; 
 constant STA_DIR : std_logic_vector (7 downto 0) :=x"ae"; 
 constant STB_DIR : std_logic_vector (7 downto 0) :=x"28"; 
 constant ADD_AB  : std_logic_vector (7 downto 0) :=x"b1"; 
 constant SUB_AB  : std_logic_vector (7 downto 0) :=x"25"; 
 constant INC_A   : std_logic_vector (7 downto 0) :=x"2b"; 
 constant DEC_A   : std_logic_vector (7 downto 0) :=x"7d"; 
 constant INC_B   : std_logic_vector (7 downto 0) :=x"b0"; 
 constant DEC_B   : std_logic_vector (7 downto 0) :=x"d3"; 
 constant AND_AB  : std_logic_vector (7 downto 0) :=x"26"; 
 constant ORR_AB  : std_logic_vector (7 downto 0) :=x"95"; 
 constant BRA     : std_logic_vector (7 downto 0) :=x"8a"; 
 constant BMI     : std_logic_vector (7 downto 0) :=x"58"; 
 constant BEQ     : std_logic_vector (7 downto 0) :=x"c7"; 
 constant BCS     : std_logic_vector (7 downto 0) :=x"1c"; 
 constant BVS     : std_logic_vector (7 downto 0) :=x"3b"; 
 constant PSH_A   : std_logic_vector (7 downto 0) :=x"7b"; 
 constant PSH_B   : std_logic_vector (7 downto 0) :=x"84"; 
 constant PSH_PC  : std_logic_vector (7 downto 0) :=x"5c"; 
 constant PLL_A   : std_logic_vector (7 downto 0) :=x"c3"; 
 constant PLL_B   : std_logic_vector (7 downto 0) :=x"47"; 
 constant PLL_PC  : std_logic_vector (7 downto 0) :=x"99"; 
 constant RTI     : std_logic_vector (7 downto 0) :=x"4b"; 
 constant STI     : std_logic_vector (7 downto 0) :=x"4a"; 
 constant add     : std_logic_vector (2 downto 0) :="000"; 
 constant sub     : std_logic_vector (2 downto 0) :="001"; 
 constant andab   : std_logic_vector (2 downto 0) :="010"; 
 constant orrab   : std_logic_vector (2 downto 0) :="011"; 
 constant inca    : std_logic_vector (2 downto 0) :="100"; 
 constant deca    : std_logic_vector (2 downto 0) :="101"; 
 constant incb    : std_logic_vector (2 downto 0) :="110"; 
 constant decb    : std_logic_vector (2 downto 0) :="111"; 
 end package instructions_core_3;