library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 
package instructions_core_1 is 
 constant LDA_IMM : std_logic_vector (7 downto 0) :=x"9b"; 
 constant LDB_IMM : std_logic_vector (7 downto 0) :=x"cf"; 
 constant LDA_DIR : std_logic_vector (7 downto 0) :=x"7a"; 
 constant LDB_DIR : std_logic_vector (7 downto 0) :=x"7d"; 
 constant STA_DIR : std_logic_vector (7 downto 0) :=x"bf"; 
 constant STB_DIR : std_logic_vector (7 downto 0) :=x"dd"; 
 constant ADD_AB  : std_logic_vector (7 downto 0) :=x"33"; 
 constant SUB_AB  : std_logic_vector (7 downto 0) :=x"74"; 
 constant INC_A   : std_logic_vector (7 downto 0) :=x"2b"; 
 constant DEC_A   : std_logic_vector (7 downto 0) :=x"c7"; 
 constant INC_B   : std_logic_vector (7 downto 0) :=x"7b"; 
 constant DEC_B   : std_logic_vector (7 downto 0) :=x"3b"; 
 constant AND_AB  : std_logic_vector (7 downto 0) :=x"93"; 
 constant ORR_AB  : std_logic_vector (7 downto 0) :=x"a6"; 
 constant BRA     : std_logic_vector (7 downto 0) :=x"ab"; 
 constant BMI     : std_logic_vector (7 downto 0) :=x"6d"; 
 constant BEQ     : std_logic_vector (7 downto 0) :=x"60"; 
 constant BCS     : std_logic_vector (7 downto 0) :=x"31"; 
 constant BVS     : std_logic_vector (7 downto 0) :=x"70"; 
 constant PSH_A   : std_logic_vector (7 downto 0) :=x"94"; 
 constant PSH_B   : std_logic_vector (7 downto 0) :=x"46"; 
 constant PSH_PC  : std_logic_vector (7 downto 0) :=x"51"; 
 constant PLL_A   : std_logic_vector (7 downto 0) :=x"8e"; 
 constant PLL_B   : std_logic_vector (7 downto 0) :=x"98"; 
 constant PLL_PC  : std_logic_vector (7 downto 0) :=x"49"; 
 constant RTI     : std_logic_vector (7 downto 0) :=x"a8"; 
 constant STI     : std_logic_vector (7 downto 0) :=x"c9"; 
 constant add     : std_logic_vector (2 downto 0) :="000"; 
 constant sub     : std_logic_vector (2 downto 0) :="001"; 
 constant andab   : std_logic_vector (2 downto 0) :="010"; 
 constant orrab   : std_logic_vector (2 downto 0) :="011"; 
 constant inca    : std_logic_vector (2 downto 0) :="100"; 
 constant deca    : std_logic_vector (2 downto 0) :="101"; 
 constant incb    : std_logic_vector (2 downto 0) :="110"; 
 constant decb    : std_logic_vector (2 downto 0) :="111"; 
 end package instructions_core_1;