library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 
package instructions_core_2 is 
 constant LDA_IMM : std_logic_vector (7 downto 0) :=x"cc"; 
 constant LDB_IMM : std_logic_vector (7 downto 0) :=x"18"; 
 constant LDA_DIR : std_logic_vector (7 downto 0) :=x"ca"; 
 constant LDB_DIR : std_logic_vector (7 downto 0) :=x"d4"; 
 constant STA_DIR : std_logic_vector (7 downto 0) :=x"32"; 
 constant STB_DIR : std_logic_vector (7 downto 0) :=x"61"; 
 constant ADD_AB  : std_logic_vector (7 downto 0) :=x"a7"; 
 constant SUB_AB  : std_logic_vector (7 downto 0) :=x"c9"; 
 constant INC_A   : std_logic_vector (7 downto 0) :=x"bb"; 
 constant DEC_A   : std_logic_vector (7 downto 0) :=x"75"; 
 constant INC_B   : std_logic_vector (7 downto 0) :=x"81"; 
 constant DEC_B   : std_logic_vector (7 downto 0) :=x"c7"; 
 constant AND_AB  : std_logic_vector (7 downto 0) :=x"1e"; 
 constant ORR_AB  : std_logic_vector (7 downto 0) :=x"aa"; 
 constant BRA     : std_logic_vector (7 downto 0) :=x"5d"; 
 constant BMI     : std_logic_vector (7 downto 0) :=x"67"; 
 constant BEQ     : std_logic_vector (7 downto 0) :=x"59"; 
 constant BCS     : std_logic_vector (7 downto 0) :=x"8b"; 
 constant BVS     : std_logic_vector (7 downto 0) :=x"b9"; 
 constant PSH_A   : std_logic_vector (7 downto 0) :=x"d7"; 
 constant PSH_B   : std_logic_vector (7 downto 0) :=x"3b"; 
 constant PSH_PC  : std_logic_vector (7 downto 0) :=x"65"; 
 constant PLL_A   : std_logic_vector (7 downto 0) :=x"4e"; 
 constant PLL_B   : std_logic_vector (7 downto 0) :=x"52"; 
 constant PLL_PC  : std_logic_vector (7 downto 0) :=x"39"; 
 constant RTI     : std_logic_vector (7 downto 0) :=x"b2"; 
 constant STI     : std_logic_vector (7 downto 0) :=x"ab"; 
 constant add     : std_logic_vector (2 downto 0) :="000"; 
 constant sub     : std_logic_vector (2 downto 0) :="001"; 
 constant andab   : std_logic_vector (2 downto 0) :="010"; 
 constant orrab   : std_logic_vector (2 downto 0) :="011"; 
 constant inca    : std_logic_vector (2 downto 0) :="100"; 
 constant deca    : std_logic_vector (2 downto 0) :="101"; 
 constant incb    : std_logic_vector (2 downto 0) :="110"; 
 constant decb    : std_logic_vector (2 downto 0) :="111"; 
 end package instructions_core_2;