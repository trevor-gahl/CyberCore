library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity char_decoder is
  port (
    char_in     : in  std_logic_vector(3 downto 0);
    led_display : out std_logic_vector(6 downto 0)
    );
end char_decoder;

architecture Behavioral of char_decoder is
begin

  decoder : process(char_in)
  begin
    case char_in is
      when "0000" =>
        led_display <= "0000001";       -- 0
      when "0001" =>
        led_display <= "1001111";       -- 1
      when "0010" =>
        led_display <= "0010010";       -- 2
      when "0011" =>
        led_display <= "0000110";       -- 3
      when "0100" =>
        led_display <= "1001100";       -- 4
      when "0101" =>
        led_display <= "0100100";       -- 5
      when "0110" =>
        led_display <= "0100000";       -- 6
      when "0111" =>
        led_display <= "0001111";       -- 7
      when "1000" =>
        led_display <= "0000000";       -- 8
      when "1001" =>
        led_display <= "0000100";       -- 9
      when "1010" =>
        led_display <= "0000010";       -- a
      when "1011" =>
        led_display <= "1100000";       -- b
      when "1100" =>
        led_display <= "0110001";       -- C
      when "1101" =>
        led_display <= "1000010";       -- d
      when "1110" =>
        led_display <= "0110000";       -- E
      when "1111" =>
        led_display <= "0111000";       -- F
      when others =>
        led_display <= "0000001";       -- 0
    end case;
  end process;

end Behavioral;
